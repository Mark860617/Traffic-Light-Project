/*LIST YOUR ULTIMATE SWAGGER IDEAS HERE
- PEDESTRIAN CROSS BUTTON
- MANUAL CONTROL VS AUTOMATION
- SHOW STATUS ON VGA
*/


module traffic_light(input [16:0] SW, input CLOCK_50, output [11:0] GPIO, input [6:0]LEDR);
	// The top level design for the traffic light intersection
	//Create wires for the slowed down clock signal and the timer.
	wire new_clock;
	wire timer;
	// Slow down the clock signal from 50 Mhz to about 1 hz
	clock_slower(.clock(CLOCK_50), .select_time(timer), .led(new_clock));
	// Adjust the different lengths before transitions of each light. 
	traffic_light_timer(.clock(new_clock), .resetn(SW[1]), .change(SW[2]), .timer(timer));
	// Output the desired signal through the GPIO pins into the indicated LEDs
	traffic_light_output(.clock(new_clock), .clock2(CLOCK_50), .resetn(SW[1]), .change(SW[2]), .set1(GPIO[4:0]), .set2(GPIO[10:5]));
endmodule

module flashLED(input clock, output reg led);
	// The module for flashing the indicated LEDs
	// Set the timer to countdown from CLOCK_50
	reg [32:0] timer = 32'd30000000;
	
	// On positive clock edge
	always @(posedge clock)
	begin
		// When the timer count is not zero decrement by 1
		if (timer != 32'd0) 
			timer <= timer - 1;
		// If timer count reaches zero, reverse LED state and reset the timer.
		else begin
			led <= ~led;
			timer <= 32'd30000000;
		end
	end
endmodule


module clock_slower(input clock, input select_time, output reg led);
	// The module for slowing down CLOCK_50's clock speed
	// Create registers for the desired countdown and the timer.
	reg [32:0] d;
	reg [32:0] timer;
	// On positive clock edge
	always @ (posedge clock)
		begin
		case (select_time)
			// Allocate the desired countdown interval depending on the select_time signal
			1'b0: d = 32'd180000000;
			1'b1: d = 32'd30000000;
			default: d = 0;
		endcase
		
		// Set timer to the desired countdown interval
		timer <= d;
		
		// When the timer count is not zero decrement timer by 1
		if (timer != 32'd0) 
			timer <= timer - 1;
		// If t1'b1imer count reaches zero, reverse LED signal and set timer to desired countdown
		else begin
			led <= ~led;
			timer <= d; // 30000000
		end
	end
endmodule


module traffic_light_timer(input clock, input resetn, input change, output reg timer);
// This is the light module for assigning the proper signals to the proper output
wire [3:0] state_sig;
control(.clock(clock), .resetn(resetn), .change(change), .out(state_sig));

 // set1 is LEDR
// set2 is LEDG
	//send signal to the breadboard
	//set1[1:0] P1 (Pedestrian Light Set 1)
	//set1[4:2] T1 (Traffic Light Set 1)
	//set2[1:0] P2 (Pedestrian Light Set 2)
	//set2[4:2] T2 (Traffic Light Set 2)
always @(*)
begin: on_off
	case(state_sig)
		4'b0000: begin //T1 R T2 G 10 secs
			timer = 1'b0;
			end
		4'b0001: begin //T1 R T2 G 10 secs
			timer = 1'b0;
			end
		4'b0010: begin //T1 R T2 Y 3 secs
			timer = 1'b1;
			end

		4'b0011: begin //T1 G T2 R 10 secs
			timer = 1'b0;
			end

		4'b0100: begin //T1 G T2 R 10 secs
			timer = 1'b0;
			end

		4'b0101: begin //T1 Y T2 R 3 secs
			timer = 1'b1;
			end
	endcase
end
endmodule



module traffic_light_output(input clock, input clock2, input resetn, input change, output reg [5:0] set1, output reg [5:0] set2);
// This is the light module for assigning the proper signals to the proper output ***LED FOR TESTING ATM***
wire [3:0] state_sig;
control(.clock(clock), .resetn(resetn), .change(change), .out(state_sig));

 // set1 is LEDR
// set2 is LEDG
	//send signal to the breadboard
	//set1[1:0] P1
	//set1[4:2] T1
	//set2[1:0] P2
	//set2[4:2] T2
wire flash_ped;
flashLED(.clock(clock2), .led(flash_ped));
always @(*)
begin: on_off
	case(state_sig)
		4'b0000: begin
			// Assign T1 to be red
			set1[4] = 1'b1;
			 set1[3] = 1'b0;
			 set1[2] = 1'b0;
			// Assign T2 to be green
			 set2[4] = 1'b0;
			 set2[3] = 1'b0;
			 set2[2] = 1'b1;
			// Assign P1 to be red
			 set1[1] = 1'b1;
			 set1[0] = 1'b0;
			// Assign P2 to be green 
			 set2[1] = 1'b0;
			 set2[0] = 1'b1;
			end
		4'b0001: begin
			// Assign T1 to be red
			 set1[4] = 1'b1;
			 set1[3] = 1'b0;
			 set1[2] = 1'b0;
			// Assign T2 to be green
			 set2[4] = 1'b0;
			 set2[3] = 1'b0;
			 set2[2] = 1'b1;
			// Assign P1 to be red
			 set1[1] = 1'b1;
			 set1[0] = 1'b0;
			 // Assign P2 to be green 
			 //Fashinf ped light on P2
			 set2[1] = flash_ped;
			 set2[0] = 1'b0;
			// 
			end
		4'b0010: begin
			// Assign T1 to be red
			 set1[4] = 1'b1;
			 set1[3] = 1'b0;
			 set1[2] = 1'b0;
			// Assign T2 to be Yellow
			 set2[4] = 1'b0;
			 set2[3] = 1'b1;
			 set2[2] = 1'b0;
			// Assign P1 to be red
			 set1[1] = 1'b1;
			 set1[0] = 1'b0;
			// Assign P2 to be Red
			 set2[1] = 1'b1;
			 set2[0] = 1'b0;
			end

		4'b0011: begin
			// Assign T1 to be green
			 set1[4] = 1'b0;
			 set1[3] = 1'b0;
			 set1[2] = 1'b1;
			// Assign T2 to be red
			 set2[4] = 1'b1;
			 set2[3] = 1'b0;
			 set2[2] = 1'b0;
			// Assign P1 to be green
			 set1[1] = 1'b0;
			 set1[0] = 1'b1;
			// Assign P2 to be red 
			 set2[1] = 1'b1;
			 set2[0] = 1'b0;
			end

		4'b0100: begin
			// Assign T1 to be green
			 set1[4] = 1'b0;
			 set1[3] = 1'b0;
			 set1[2] = 1'b1;
			// Assign T2 to be red
			 set2[4] = 1'b1;
			 set2[3] = 1'b0;
			 set2[2] = 1'b0;
			// Assign P1 to be green
			 set1[1] = flash_ped;
			 set1[0] = 1'b0;
			// Assign P2 to be red 
			 set2[1] = 1'b1;
			 set2[0] = 1'b0;
			end

		4'b0101: begin
			// Assign T1 to be yellow
			 set1[4] = 1'b0;
			 set1[3] = 1'b1;
			 set1[2] = 1'b0;
			// Assign T2 to be red
			 set2[4] = 1'b1;
			 set2[3] = 1'b0;
			 set2[2] = 1'b0;
			//Assign P1 to be red
			 set1[1] = 1'b1;
			 set1[0] = 1'b0;
			// Assign P2 to be red 
			 set2[1] = 1'b1;
			 set2[0] = 1'b0;
			end
	endcase
end
endmodule



module control(input clock, input resetn, input change, output [3:0] out);
	// The fsm to determine the state of the traffic/pedestrian lights
	reg [3:0] curr, next;

	//State A is T1 red, T2 green, p1 red, p2 green
	localparam A = 4'b0000, B = 4'b0001, C = 4'b0010, D = 4'b0011, E = 4'b0100, F = 4'b0101;

	always @(*)
	begin: state_table
		case(curr)
			A: begin
				if (!change) next <= A;
				else next <= B;
			end
			B: begin
				if (!change) next <= B;
				else next <= C;	
			end
			C: begin
				if (!change) next <= C;
				else next <= D;	
			end
			D: begin
				if (!change) next <= D;
				else next <= E;	
			end
			E: begin
				if (!change) next <= E;
				else next <= F;	
			end
			F: begin
				if (!change) next <= F;
				else next <= A;	
			end
			default: next <= A;
		endcase
	end

	always @(posedge clock)
		begin: flip_flops
			if (resetn == 1'b0)
				curr <= A;
			else
				curr <= next;
		end

	assign out = curr;

endmodule

module hex_decoder(hex_digit, segments);
    input hex_digit; // change it back to [3:0]
    output reg [6:0] segments;

    always @(*)
        case (hex_digit)
            4'h0: segments = 7'b100_0000;
            4'h1: segments = 7'b111_1001;
            4'h2: segments = 7'b010_0100;
            4'h3: segments = 7'b011_0000;
            4'h4: segments = 7'b001_1001;
            4'h5: segments = 7'b001_0010;
            4'h6: segments = 7'b000_0010;
            4'h7: segments = 7'b111_1000;
            4'h8: segments = 7'b000_0000;
            4'h9: segments = 7'b001_1000;
            4'hA: segments = 7'b000_1000;
            4'hB: segments = 7'b000_0011;
            4'hC: segments = 7'b100_0110;
            4'hD: segments = 7'b010_0001;
            4'hE: segments = 7'b000_0110;
            4'hF: segments = 7'b000_1110;
            default: segments = 7'h7f;
        endcase
endmodule

